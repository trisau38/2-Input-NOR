.title nor_2_inp
.include techfile130.txt

vdd vdd 0 1.2

vA A 0 PULSE(0 1.2 2NS 2NS 2NS 50NS 100NS)
vB B 0 PULSE(0 1.2 20NS 2NS 2NS 50NS 100NS)

Mp1 1 A vdd vdd pmos l=120n w=2880n
Mp2 vout B 1 vdd pmos l=120n w=2880n

Mn1 vout A 0 0 nmos l=120n w=480n
Mn2 vout B 0 0 nmos l=120n w=480n


.tran 0.1n 200n 0 0.1n

.control
run 
plot v(A) v(B) v(vout)
.endc
.end
